`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04.10.2022 08:44:29
// Design Name: 
// Module Name: mux_in_time_4x4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux_in_time_4x4(
    input [4:0] dato0,
    input [4:0] dato1,
    input [4:0] dato2,
    input [4:0] dato3,
    input clk,
    output [3:0] segm,
    output [3:0] transistor
    );
endmodule
