`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04.10.2022 08:41:39
// Design Name: 
// Module Name: adder_subs
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module adder_subs(
    input [3:0] a,
    input [3:0] b,
    input sum_rest,
    input clk,
    output [6:0] segm,
    output [3:0] transistor
    );
endmodule
